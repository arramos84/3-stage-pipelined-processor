module app(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h27bdffa8;
30'h00000001: inst = 32'hafbf0050;
30'h00000002: inst = 32'hafb00040;
30'h00000003: inst = 32'hafb10044;
30'h00000004: inst = 32'hafb20048;
30'h00000005: inst = 32'h3c021fff;
30'h00000006: inst = 32'h34430000;
30'h00000007: inst = 32'hafa00020;
30'h00000008: inst = 32'h34440004;
30'h00000009: inst = 32'hac600000;
30'h0000000a: inst = 32'h34430010;
30'h0000000b: inst = 32'hac800000;
30'h0000000c: inst = 32'h34440014;
30'h0000000d: inst = 32'hac600000;
30'h0000000e: inst = 32'h34430008;
30'h0000000f: inst = 32'hac800000;
30'h00000010: inst = 32'h24040001;
30'h00000011: inst = 32'h34420018;
30'h00000012: inst = 32'hac600000;
30'h00000013: inst = 32'hac440000;
30'h00000014: inst = 32'h40804800;
30'h00000015: inst = 32'h00000000;
30'h00000016: inst = 32'h341a8c01;
30'h00000017: inst = 32'h00000000;
30'h00000018: inst = 32'h409a6000;
30'h00000019: inst = 32'h00000000;
30'h0000001a: inst = 32'h3c021fff;
30'h0000001b: inst = 32'h34420008;
30'h0000001c: inst = 32'h8c420000;
30'h0000001d: inst = 32'h00000000;
30'h0000001e: inst = 32'h24030071;
30'h0000001f: inst = 32'h0062182a;
30'h00000020: inst = 32'h14600023;
30'h00000021: inst = 32'h00000000;
30'h00000022: inst = 32'h24030052;
30'h00000023: inst = 32'h10430055;
30'h00000024: inst = 32'h00000000;
30'h00000025: inst = 32'h24030056;
30'h00000026: inst = 32'h1443fff3;
30'h00000027: inst = 32'h00000000;
30'h00000028: inst = 32'h3c021fff;
30'h00000029: inst = 32'h34430010;
30'h0000002a: inst = 32'h8c640000;
30'h0000002b: inst = 32'h00000000;
30'h0000002c: inst = 32'h2405003c;
30'h0000002d: inst = 32'h34500014;
30'h0000002e: inst = 32'h0c0000c0;
30'h0000002f: inst = 32'h00000000;
30'h00000030: inst = 32'h8e030000;
30'h00000031: inst = 32'h00000000;
30'h00000032: inst = 32'h00431021;
30'h00000033: inst = 32'hafa20024;
30'h00000034: inst = 32'hafa0003c;
30'h00000035: inst = 32'h3c0205f5;
30'h00000036: inst = 32'h3442e0ff;
30'h00000037: inst = 32'h8fa3003c;
30'h00000038: inst = 32'h00000000;
30'h00000039: inst = 32'h0043102b;
30'h0000003a: inst = 32'h1440006b;
30'h0000003b: inst = 32'h00000000;
30'h0000003c: inst = 32'h0c000243;
30'h0000003d: inst = 32'h00000000;
30'h0000003e: inst = 32'h8fa2003c;
30'h0000003f: inst = 32'h00000000;
30'h00000040: inst = 32'h24420001;
30'h00000041: inst = 32'hafa2003c;
30'h00000042: inst = 32'h08000035;
30'h00000043: inst = 32'h00000000;
30'h00000044: inst = 32'h24030076;
30'h00000045: inst = 32'h1043004f;
30'h00000046: inst = 32'h00000000;
30'h00000047: inst = 32'h24030072;
30'h00000048: inst = 32'h1443ffd1;
30'h00000049: inst = 32'h00000000;
30'h0000004a: inst = 32'h3c021fff;
30'h0000004b: inst = 32'h34500010;
30'h0000004c: inst = 32'h8e040000;
30'h0000004d: inst = 32'h00000000;
30'h0000004e: inst = 32'h2411003c;
30'h0000004f: inst = 32'h34520014;
30'h00000050: inst = 32'h00112821;
30'h00000051: inst = 32'h0c0000c0;
30'h00000052: inst = 32'h00000000;
30'h00000053: inst = 32'h8e430000;
30'h00000054: inst = 32'h00000000;
30'h00000055: inst = 32'h00431021;
30'h00000056: inst = 32'hafa20024;
30'h00000057: inst = 32'h0c000212;
30'h00000058: inst = 32'h00000000;
30'h00000059: inst = 32'h8e040000;
30'h0000005a: inst = 32'h00000000;
30'h0000005b: inst = 32'h00112821;
30'h0000005c: inst = 32'h0c0000c0;
30'h0000005d: inst = 32'h00000000;
30'h0000005e: inst = 32'h8e430000;
30'h0000005f: inst = 32'h00000000;
30'h00000060: inst = 32'h00431021;
30'h00000061: inst = 32'hafa20028;
30'h00000062: inst = 32'h8fa30024;
30'h00000063: inst = 32'h00000000;
30'h00000064: inst = 32'h00432023;
30'h00000065: inst = 32'hafa4002c;
30'h00000066: inst = 32'h00112821;
30'h00000067: inst = 32'h0c0000dd;
30'h00000068: inst = 32'h00000000;
30'h00000069: inst = 32'hafa20030;
30'h0000006a: inst = 32'h8fa4002c;
30'h0000006b: inst = 32'h00000000;
30'h0000006c: inst = 32'h00112821;
30'h0000006d: inst = 32'h0c0000fb;
30'h0000006e: inst = 32'h00000000;
30'h0000006f: inst = 32'hafa20034;
30'h00000070: inst = 32'h8fa40030;
30'h00000071: inst = 32'h00000000;
30'h00000072: inst = 32'h00022821;
30'h00000073: inst = 32'h0c000114;
30'h00000074: inst = 32'h00000000;
30'h00000075: inst = 32'h0c000162;
30'h00000076: inst = 32'h00000000;
30'h00000077: inst = 32'h0800001a;
30'h00000078: inst = 32'h00000000;
30'h00000079: inst = 32'h3c021fff;
30'h0000007a: inst = 32'h34430010;
30'h0000007b: inst = 32'h8c640000;
30'h0000007c: inst = 32'h00000000;
30'h0000007d: inst = 32'h2405003c;
30'h0000007e: inst = 32'h34500014;
30'h0000007f: inst = 32'h0c0000c0;
30'h00000080: inst = 32'h00000000;
30'h00000081: inst = 32'h8e030000;
30'h00000082: inst = 32'h00000000;
30'h00000083: inst = 32'h00431021;
30'h00000084: inst = 32'hafa20024;
30'h00000085: inst = 32'hafa00038;
30'h00000086: inst = 32'h3c0205f5;
30'h00000087: inst = 32'h3442e0ff;
30'h00000088: inst = 32'h8fa30038;
30'h00000089: inst = 32'h00000000;
30'h0000008a: inst = 32'h0043102b;
30'h0000008b: inst = 32'h1440001a;
30'h0000008c: inst = 32'h00000000;
30'h0000008d: inst = 32'h0c000224;
30'h0000008e: inst = 32'h00000000;
30'h0000008f: inst = 32'h8fa20038;
30'h00000090: inst = 32'h00000000;
30'h00000091: inst = 32'h24420001;
30'h00000092: inst = 32'hafa20038;
30'h00000093: inst = 32'h08000086;
30'h00000094: inst = 32'h00000000;
30'h00000095: inst = 32'h3c021fff;
30'h00000096: inst = 32'h34500010;
30'h00000097: inst = 32'h8e040000;
30'h00000098: inst = 32'h00000000;
30'h00000099: inst = 32'h2411003c;
30'h0000009a: inst = 32'h34520014;
30'h0000009b: inst = 32'h00112821;
30'h0000009c: inst = 32'h0c0000c0;
30'h0000009d: inst = 32'h00000000;
30'h0000009e: inst = 32'h8e430000;
30'h0000009f: inst = 32'h00000000;
30'h000000a0: inst = 32'h00431021;
30'h000000a1: inst = 32'hafa20024;
30'h000000a2: inst = 32'h0c00022b;
30'h000000a3: inst = 32'h00000000;
30'h000000a4: inst = 32'h08000059;
30'h000000a5: inst = 32'h00000000;
30'h000000a6: inst = 32'h3c021fff;
30'h000000a7: inst = 32'h34430010;
30'h000000a8: inst = 32'h8c640000;
30'h000000a9: inst = 32'h00000000;
30'h000000aa: inst = 32'h2410003c;
30'h000000ab: inst = 32'h34510014;
30'h000000ac: inst = 32'h00102821;
30'h000000ad: inst = 32'h0c0000c0;
30'h000000ae: inst = 32'h00000000;
30'h000000af: inst = 32'h8e230000;
30'h000000b0: inst = 32'h00000000;
30'h000000b1: inst = 32'h00431021;
30'h000000b2: inst = 32'hafa20028;
30'h000000b3: inst = 32'h8fa30024;
30'h000000b4: inst = 32'h00000000;
30'h000000b5: inst = 32'h00432023;
30'h000000b6: inst = 32'hafa4002c;
30'h000000b7: inst = 32'h00102821;
30'h000000b8: inst = 32'h0c0000dd;
30'h000000b9: inst = 32'h00000000;
30'h000000ba: inst = 32'hafa20030;
30'h000000bb: inst = 32'h8fa4002c;
30'h000000bc: inst = 32'h00000000;
30'h000000bd: inst = 32'h00102821;
30'h000000be: inst = 32'h0800006d;
30'h000000bf: inst = 32'h00000000;
30'h000000c0: inst = 32'h27bdffe0;
30'h000000c1: inst = 32'hafa40010;
30'h000000c2: inst = 32'hafa50014;
30'h000000c3: inst = 32'hafa00018;
30'h000000c4: inst = 32'hafa0001c;
30'h000000c5: inst = 32'h8fa2001c;
30'h000000c6: inst = 32'h00000000;
30'h000000c7: inst = 32'h8fa30014;
30'h000000c8: inst = 32'h00000000;
30'h000000c9: inst = 32'h0043102a;
30'h000000ca: inst = 32'h1040000d;
30'h000000cb: inst = 32'h00000000;
30'h000000cc: inst = 32'h8fa20010;
30'h000000cd: inst = 32'h00000000;
30'h000000ce: inst = 32'h8fa30018;
30'h000000cf: inst = 32'h00000000;
30'h000000d0: inst = 32'h00621021;
30'h000000d1: inst = 32'hafa20018;
30'h000000d2: inst = 32'h8fa2001c;
30'h000000d3: inst = 32'h00000000;
30'h000000d4: inst = 32'h24420001;
30'h000000d5: inst = 32'hafa2001c;
30'h000000d6: inst = 32'h080000c5;
30'h000000d7: inst = 32'h00000000;
30'h000000d8: inst = 32'h8fa20018;
30'h000000d9: inst = 32'h00000000;
30'h000000da: inst = 32'h27bd0020;
30'h000000db: inst = 32'h03e00008;
30'h000000dc: inst = 32'h00000000;
30'h000000dd: inst = 32'h27bdffe0;
30'h000000de: inst = 32'hafa40010;
30'h000000df: inst = 32'hafa50014;
30'h000000e0: inst = 32'hafa00018;
30'h000000e1: inst = 32'h8fa20010;
30'h000000e2: inst = 32'h00000000;
30'h000000e3: inst = 32'hafa2001c;
30'h000000e4: inst = 32'h8fa2001c;
30'h000000e5: inst = 32'h00000000;
30'h000000e6: inst = 32'h8fa30014;
30'h000000e7: inst = 32'h00000000;
30'h000000e8: inst = 32'h0043102a;
30'h000000e9: inst = 32'h1440000c;
30'h000000ea: inst = 32'h00000000;
30'h000000eb: inst = 32'h8fa20018;
30'h000000ec: inst = 32'h00000000;
30'h000000ed: inst = 32'h24420001;
30'h000000ee: inst = 32'hafa20018;
30'h000000ef: inst = 32'h8fa20014;
30'h000000f0: inst = 32'h00000000;
30'h000000f1: inst = 32'h8fa3001c;
30'h000000f2: inst = 32'h00000000;
30'h000000f3: inst = 32'h00621023;
30'h000000f4: inst = 32'h080000e3;
30'h000000f5: inst = 32'h00000000;
30'h000000f6: inst = 32'h8fa20018;
30'h000000f7: inst = 32'h00000000;
30'h000000f8: inst = 32'h27bd0020;
30'h000000f9: inst = 32'h03e00008;
30'h000000fa: inst = 32'h00000000;
30'h000000fb: inst = 32'h27bdffe0;
30'h000000fc: inst = 32'hafa40010;
30'h000000fd: inst = 32'hafa50014;
30'h000000fe: inst = 32'h8fa20010;
30'h000000ff: inst = 32'h00000000;
30'h00000100: inst = 32'hafa20018;
30'h00000101: inst = 32'h8fa20018;
30'h00000102: inst = 32'h00000000;
30'h00000103: inst = 32'h8fa30014;
30'h00000104: inst = 32'h00000000;
30'h00000105: inst = 32'h0043102a;
30'h00000106: inst = 32'h14400008;
30'h00000107: inst = 32'h00000000;
30'h00000108: inst = 32'h8fa20014;
30'h00000109: inst = 32'h00000000;
30'h0000010a: inst = 32'h8fa30018;
30'h0000010b: inst = 32'h00000000;
30'h0000010c: inst = 32'h00621023;
30'h0000010d: inst = 32'h08000100;
30'h0000010e: inst = 32'h00000000;
30'h0000010f: inst = 32'h8fa20018;
30'h00000110: inst = 32'h00000000;
30'h00000111: inst = 32'h27bd0020;
30'h00000112: inst = 32'h03e00008;
30'h00000113: inst = 32'h00000000;
30'h00000114: inst = 32'h27bdffb8;
30'h00000115: inst = 32'hafbf0040;
30'h00000116: inst = 32'hafb00038;
30'h00000117: inst = 32'hafa40020;
30'h00000118: inst = 32'hafa50024;
30'h00000119: inst = 32'hafa0002c;
30'h0000011a: inst = 32'h8fa20020;
30'h0000011b: inst = 32'h00000000;
30'h0000011c: inst = 32'hafa20028;
30'h0000011d: inst = 32'hafa00034;
30'h0000011e: inst = 32'h8fa20024;
30'h0000011f: inst = 32'h00000000;
30'h00000120: inst = 32'hafa20030;
30'h00000121: inst = 32'h8fa20028;
30'h00000122: inst = 32'h00000000;
30'h00000123: inst = 32'h2842000a;
30'h00000124: inst = 32'h1440000b;
30'h00000125: inst = 32'h00000000;
30'h00000126: inst = 32'h8fa20028;
30'h00000127: inst = 32'h00000000;
30'h00000128: inst = 32'h2442fff6;
30'h00000129: inst = 32'hafa20028;
30'h0000012a: inst = 32'h8fa2002c;
30'h0000012b: inst = 32'h00000000;
30'h0000012c: inst = 32'h24420001;
30'h0000012d: inst = 32'hafa2002c;
30'h0000012e: inst = 32'h08000121;
30'h0000012f: inst = 32'h00000000;
30'h00000130: inst = 32'h8fa4002c;
30'h00000131: inst = 32'h00000000;
30'h00000132: inst = 32'h3c101000;
30'h00000133: inst = 32'h0c0001df;
30'h00000134: inst = 32'h00000000;
30'h00000135: inst = 32'h26030974;
30'h00000136: inst = 32'ha0620000;
30'h00000137: inst = 32'h8fa40028;
30'h00000138: inst = 32'h00000000;
30'h00000139: inst = 32'h3c101000;
30'h0000013a: inst = 32'h0c0001df;
30'h0000013b: inst = 32'h00000000;
30'h0000013c: inst = 32'h26030978;
30'h0000013d: inst = 32'ha0620000;
30'h0000013e: inst = 32'h8fa20030;
30'h0000013f: inst = 32'h00000000;
30'h00000140: inst = 32'h2842000a;
30'h00000141: inst = 32'h1440000b;
30'h00000142: inst = 32'h00000000;
30'h00000143: inst = 32'h8fa20030;
30'h00000144: inst = 32'h00000000;
30'h00000145: inst = 32'h2442fff6;
30'h00000146: inst = 32'hafa20030;
30'h00000147: inst = 32'h8fa20034;
30'h00000148: inst = 32'h00000000;
30'h00000149: inst = 32'h24420001;
30'h0000014a: inst = 32'hafa20034;
30'h0000014b: inst = 32'h0800013e;
30'h0000014c: inst = 32'h00000000;
30'h0000014d: inst = 32'h8fa40034;
30'h0000014e: inst = 32'h00000000;
30'h0000014f: inst = 32'h3c101000;
30'h00000150: inst = 32'h0c0001df;
30'h00000151: inst = 32'h00000000;
30'h00000152: inst = 32'h2603097c;
30'h00000153: inst = 32'ha0620000;
30'h00000154: inst = 32'h8fa40030;
30'h00000155: inst = 32'h00000000;
30'h00000156: inst = 32'h3c101000;
30'h00000157: inst = 32'h0c0001df;
30'h00000158: inst = 32'h00000000;
30'h00000159: inst = 32'h26030970;
30'h0000015a: inst = 32'ha0620000;
30'h0000015b: inst = 32'h8fb00038;
30'h0000015c: inst = 32'h00000000;
30'h0000015d: inst = 32'h8fbf0040;
30'h0000015e: inst = 32'h00000000;
30'h0000015f: inst = 32'h27bd0048;
30'h00000160: inst = 32'h03e00008;
30'h00000161: inst = 32'h00000000;
30'h00000162: inst = 32'h27bdffe8;
30'h00000163: inst = 32'h3c021000;
30'h00000164: inst = 32'h24420980;
30'h00000165: inst = 32'h2403000a;
30'h00000166: inst = 32'h24040009;
30'h00000167: inst = 32'ha0430000;
30'h00000168: inst = 32'h2405004d;
30'h00000169: inst = 32'ha0440001;
30'h0000016a: inst = 32'h2404006f;
30'h0000016b: inst = 32'ha0450002;
30'h0000016c: inst = 32'h24050064;
30'h0000016d: inst = 32'ha0440003;
30'h0000016e: inst = 32'h24040065;
30'h0000016f: inst = 32'ha0450004;
30'h00000170: inst = 32'h2405003a;
30'h00000171: inst = 32'ha0440005;
30'h00000172: inst = 32'h3c061fff;
30'h00000173: inst = 32'h24070020;
30'h00000174: inst = 32'ha0450006;
30'h00000175: inst = 32'h34c60008;
30'h00000176: inst = 32'ha0470007;
30'h00000177: inst = 32'h8cc60000;
30'h00000178: inst = 32'h00000000;
30'h00000179: inst = 32'ha0460008;
30'h0000017a: inst = 32'h24060054;
30'h0000017b: inst = 32'ha0470009;
30'h0000017c: inst = 32'h24080069;
30'h0000017d: inst = 32'ha046000a;
30'h0000017e: inst = 32'h2406006d;
30'h0000017f: inst = 32'ha048000b;
30'h00000180: inst = 32'ha046000c;
30'h00000181: inst = 32'ha044000d;
30'h00000182: inst = 32'h3c041000;
30'h00000183: inst = 32'ha045000e;
30'h00000184: inst = 32'h24840974;
30'h00000185: inst = 32'ha047000f;
30'h00000186: inst = 32'h90840000;
30'h00000187: inst = 32'h00000000;
30'h00000188: inst = 32'h3c061000;
30'h00000189: inst = 32'h24c60978;
30'h0000018a: inst = 32'ha0440010;
30'h0000018b: inst = 32'h90c40000;
30'h0000018c: inst = 32'h00000000;
30'h0000018d: inst = 32'h3c061000;
30'h0000018e: inst = 32'ha0440011;
30'h0000018f: inst = 32'h24c4097c;
30'h00000190: inst = 32'ha0450012;
30'h00000191: inst = 32'h90840000;
30'h00000192: inst = 32'h00000000;
30'h00000193: inst = 32'h3c051000;
30'h00000194: inst = 32'h24a50970;
30'h00000195: inst = 32'ha0440013;
30'h00000196: inst = 32'h90a40000;
30'h00000197: inst = 32'h00000000;
30'h00000198: inst = 32'ha0440014;
30'h00000199: inst = 32'ha0430015;
30'h0000019a: inst = 32'h24040000;
30'h0000019b: inst = 32'ha0430016;
30'h0000019c: inst = 32'h3c038000;
30'h0000019d: inst = 32'ha0440017;
30'h0000019e: inst = 32'h34620000;
30'h0000019f: inst = 32'hafa00010;
30'h000001a0: inst = 32'h8c420000;
30'h000001a1: inst = 32'h00000000;
30'h000001a2: inst = 32'h30420001;
30'h000001a3: inst = 32'h1040000f;
30'h000001a4: inst = 32'h00000000;
30'h000001a5: inst = 32'h3c021000;
30'h000001a6: inst = 32'h24420980;
30'h000001a7: inst = 32'h8fa30010;
30'h000001a8: inst = 32'h00000000;
30'h000001a9: inst = 32'h00431021;
30'h000001aa: inst = 32'h90420000;
30'h000001ab: inst = 32'h00000000;
30'h000001ac: inst = 32'h3c038000;
30'h000001ad: inst = 32'h34630008;
30'h000001ae: inst = 32'hac620000;
30'h000001af: inst = 32'h8fa20010;
30'h000001b0: inst = 32'h00000000;
30'h000001b1: inst = 32'h24420001;
30'h000001b2: inst = 32'hafa20010;
30'h000001b3: inst = 32'h3c021000;
30'h000001b4: inst = 32'h24420980;
30'h000001b5: inst = 32'h8fa30010;
30'h000001b6: inst = 32'h00000000;
30'h000001b7: inst = 32'h00431021;
30'h000001b8: inst = 32'h3c031fff;
30'h000001b9: inst = 32'h90420000;
30'h000001ba: inst = 32'h00000000;
30'h000001bb: inst = 32'h34640000;
30'h000001bc: inst = 32'h3463001c;
30'h000001bd: inst = 32'h8c840000;
30'h000001be: inst = 32'h00000000;
30'h000001bf: inst = 32'h00831821;
30'h000001c0: inst = 32'ha0620000;
30'h000001c1: inst = 32'h90620000;
30'h000001c2: inst = 32'h00000000;
30'h000001c3: inst = 32'h10400015;
30'h000001c4: inst = 32'h00000000;
30'h000001c5: inst = 32'h3c021fff;
30'h000001c6: inst = 32'h34420000;
30'h000001c7: inst = 32'h8c420000;
30'h000001c8: inst = 32'h00000000;
30'h000001c9: inst = 32'h240307ff;
30'h000001ca: inst = 32'h14430006;
30'h000001cb: inst = 32'h00000000;
30'h000001cc: inst = 32'h3c021fff;
30'h000001cd: inst = 32'h34420000;
30'h000001ce: inst = 32'hac400000;
30'h000001cf: inst = 32'h080001af;
30'h000001d0: inst = 32'h00000000;
30'h000001d1: inst = 32'h3c021fff;
30'h000001d2: inst = 32'h34420000;
30'h000001d3: inst = 32'h8c430000;
30'h000001d4: inst = 32'h00000000;
30'h000001d5: inst = 32'h24630001;
30'h000001d6: inst = 32'hac430000;
30'h000001d7: inst = 32'h080001af;
30'h000001d8: inst = 32'h00000000;
30'h000001d9: inst = 32'h3c021fff;
30'h000001da: inst = 32'h34420008;
30'h000001db: inst = 32'hac400000;
30'h000001dc: inst = 32'h27bd0018;
30'h000001dd: inst = 32'h03e00008;
30'h000001de: inst = 32'h00000000;
30'h000001df: inst = 32'h27bdffe8;
30'h000001e0: inst = 32'h24020009;
30'h000001e1: inst = 32'hafa40014;
30'h000001e2: inst = 32'h0044102b;
30'h000001e3: inst = 32'h14400027;
30'h000001e4: inst = 32'h00000000;
30'h000001e5: inst = 32'h3c021000;
30'h000001e6: inst = 32'h00041880;
30'h000001e7: inst = 32'h24420934;
30'h000001e8: inst = 32'h00621021;
30'h000001e9: inst = 32'h8c420000;
30'h000001ea: inst = 32'h00000000;
30'h000001eb: inst = 32'h00400008;
30'h000001ec: inst = 32'h00000000;
30'h000001ed: inst = 32'h24020030;
30'h000001ee: inst = 32'h0800020c;
30'h000001ef: inst = 32'h00000000;
30'h000001f0: inst = 32'h24020031;
30'h000001f1: inst = 32'h0800020c;
30'h000001f2: inst = 32'h00000000;
30'h000001f3: inst = 32'h24020032;
30'h000001f4: inst = 32'h0800020c;
30'h000001f5: inst = 32'h00000000;
30'h000001f6: inst = 32'h24020033;
30'h000001f7: inst = 32'h0800020c;
30'h000001f8: inst = 32'h00000000;
30'h000001f9: inst = 32'h24020034;
30'h000001fa: inst = 32'h0800020c;
30'h000001fb: inst = 32'h00000000;
30'h000001fc: inst = 32'h24020035;
30'h000001fd: inst = 32'h0800020c;
30'h000001fe: inst = 32'h00000000;
30'h000001ff: inst = 32'h24020036;
30'h00000200: inst = 32'h0800020c;
30'h00000201: inst = 32'h00000000;
30'h00000202: inst = 32'h24020037;
30'h00000203: inst = 32'h0800020c;
30'h00000204: inst = 32'h00000000;
30'h00000205: inst = 32'h24020038;
30'h00000206: inst = 32'h0800020c;
30'h00000207: inst = 32'h00000000;
30'h00000208: inst = 32'h24020039;
30'h00000209: inst = 32'h0800020c;
30'h0000020a: inst = 32'h00000000;
30'h0000020b: inst = 32'h24020023;
30'h0000020c: inst = 32'ha3a20010;
30'h0000020d: inst = 32'h93a20010;
30'h0000020e: inst = 32'h00000000;
30'h0000020f: inst = 32'h27bd0018;
30'h00000210: inst = 32'h03e00008;
30'h00000211: inst = 32'h00000000;
30'h00000212: inst = 32'h27bdffe8;
30'h00000213: inst = 32'hafa00010;
30'h00000214: inst = 32'h3c0205f5;
30'h00000215: inst = 32'h3442e0ff;
30'h00000216: inst = 32'h8fa30010;
30'h00000217: inst = 32'h00000000;
30'h00000218: inst = 32'h0043102a;
30'h00000219: inst = 32'h14400007;
30'h0000021a: inst = 32'h00000000;
30'h0000021b: inst = 32'h8fa20010;
30'h0000021c: inst = 32'h00000000;
30'h0000021d: inst = 32'h24420001;
30'h0000021e: inst = 32'hafa20010;
30'h0000021f: inst = 32'h08000214;
30'h00000220: inst = 32'h00000000;
30'h00000221: inst = 32'h27bd0018;
30'h00000222: inst = 32'h03e00008;
30'h00000223: inst = 32'h00000000;
30'h00000224: inst = 32'h27bdffe8;
30'h00000225: inst = 32'h24020001;
30'h00000226: inst = 32'hafa00010;
30'h00000227: inst = 32'hafa20010;
30'h00000228: inst = 32'h27bd0018;
30'h00000229: inst = 32'h03e00008;
30'h0000022a: inst = 32'h00000000;
30'h0000022b: inst = 32'h27bdfff0;
30'h0000022c: inst = 32'h3c021fff;
30'h0000022d: inst = 32'h3442000c;
30'h0000022e: inst = 32'hac400000;
30'h0000022f: inst = 32'h3c021fff;
30'h00000230: inst = 32'h3c0305f5;
30'h00000231: inst = 32'h3442000c;
30'h00000232: inst = 32'h3463e0ff;
30'h00000233: inst = 32'h8c420000;
30'h00000234: inst = 32'h00000000;
30'h00000235: inst = 32'h0062102b;
30'h00000236: inst = 32'h14400009;
30'h00000237: inst = 32'h00000000;
30'h00000238: inst = 32'h3c021fff;
30'h00000239: inst = 32'h3442000c;
30'h0000023a: inst = 32'h8c430000;
30'h0000023b: inst = 32'h00000000;
30'h0000023c: inst = 32'h24630001;
30'h0000023d: inst = 32'hac430000;
30'h0000023e: inst = 32'h0800022f;
30'h0000023f: inst = 32'h00000000;
30'h00000240: inst = 32'h27bd0010;
30'h00000241: inst = 32'h03e00008;
30'h00000242: inst = 32'h00000000;
30'h00000243: inst = 32'h27bdfff0;
30'h00000244: inst = 32'h3c021fff;
30'h00000245: inst = 32'h3442000c;
30'h00000246: inst = 32'h8c430000;
30'h00000247: inst = 32'h00000000;
30'h00000248: inst = 32'h24630001;
30'h00000249: inst = 32'hac430000;
30'h0000024a: inst = 32'h27bd0010;
30'h0000024b: inst = 32'h03e00008;
30'h0000024c: inst = 32'h00000000;
30'h0000024d: inst = 32'h100007b4;
30'h0000024e: inst = 32'h100007c0;
30'h0000024f: inst = 32'h100007cc;
30'h00000250: inst = 32'h100007d8;
30'h00000251: inst = 32'h100007e4;
30'h00000252: inst = 32'h100007f0;
30'h00000253: inst = 32'h100007fc;
30'h00000254: inst = 32'h10000808;
30'h00000255: inst = 32'h10000814;
30'h00000256: inst = 32'h10000820;
30'h00000257: inst = 32'h30313233;
30'h00000258: inst = 32'h34353637;
30'h00000259: inst = 32'h38390000;
30'h0000025a: inst = 32'h00000000;
default:      inst = 32'h00000000;
endcase
end
endmodule
