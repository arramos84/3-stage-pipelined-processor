module asmtest(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h24170000;
30'h00000001: inst = 32'h24100020;
30'h00000002: inst = 32'h24080020;
30'h00000003: inst = 32'h1510001a;
30'h00000004: inst = 32'h26f70001;
30'h00000005: inst = 32'h24100001;
30'h00000006: inst = 32'h24081000;
30'h00000007: inst = 32'h001080c0;
30'h00000008: inst = 32'h15100015;
30'h00000009: inst = 32'h26f7000a;
30'h0000000a: inst = 32'h24101000;
30'h0000000b: inst = 32'h24080001;
30'h0000000c: inst = 32'h001080c2;
30'h0000000d: inst = 32'h15100010;
30'h0000000e: inst = 32'h26f7000b;
30'h0000000f: inst = 32'h3c101111;
30'h00000010: inst = 32'h36101000;
30'h00000011: inst = 32'h3c081111;
30'h00000012: inst = 32'h35081110;
30'h00000013: inst = 32'h00108083;
30'h00000014: inst = 32'h15100009;
30'h00000015: inst = 32'h26f7000c;
30'h00000016: inst = 32'h24110003;
30'h00000017: inst = 32'h24100001;
30'h00000018: inst = 32'h24081000;
30'h00000019: inst = 32'h02308007;
30'h0000001a: inst = 32'h15100003;
30'h0000001b: inst = 32'h26f7000d;
30'h0000001c: inst = 32'h08000021;
30'h0000001d: inst = 32'h00000000;
30'h0000001e: inst = 32'h3c108000;
30'h0000001f: inst = 32'h36100008;
30'h00000020: inst = 32'hae170000;
30'h00000021: inst = 32'h241100ff;
30'h00000022: inst = 32'h3c108000;
30'h00000023: inst = 32'h36100008;
30'h00000024: inst = 32'hae110000;
default:      inst = 32'h00000000;
endcase
end
endmodule
